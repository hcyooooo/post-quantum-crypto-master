`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Technical University of Munich
// Engineer: Tim Fritzmann
// 
// Create Date: 01/27/2020
// Module Name: mul_ternary_top_tb
// Project Name: Post-Quantum Cryptography
// 
//////////////////////////////////////////////////////////////////////////////////


`define REF_CLK_PERIOD   (2*15.25us)  // 32.786 kHz --> FLL reset value --> 50 MHz
`define CLK_PERIOD       40.00ns      // 25 MHz

module mul_ternary_top_tb();
    parameter PARAM_N = 512;

    logic clk;
    logic rst;
    logic enable_write;
    logic enable_calc;
    logic enable_read;
    logic [31:0] in_1;
    logic [31:0] in_2;
    logic [31:0] out_1;
    logic ready;
    
    logic [7:0] poly_gen [PARAM_N-1:0] = {104, 139, 61, 90, 180, 237, 92, 147, 131, 144, 129, 60, 141, 242, 9, 173, 91, 175, 116, 9, 202, 203, 247, 235, 222, 229, 231, 80, 114, 155, 234, 96, 52, 68, 248, 150, 238, 234, 97, 179, 132, 39, 127, 142, 233, 110, 77, 32, 133, 8, 157, 207, 187, 131, 200, 34, 160, 140, 106, 236, 146, 69, 196, 54, 25, 153, 97, 162, 51, 175, 166, 249, 209, 79, 26, 90, 169, 201, 61, 97, 133, 99, 20, 168, 54, 82, 103, 135, 120, 26, 115, 40, 137, 63, 27, 121, 66, 14, 168, 88, 54, 108, 144, 129, 177, 96, 65, 122, 134, 59, 119, 152, 193, 84, 173, 166, 147, 92, 126, 216, 132, 49, 95, 44, 198, 25, 41, 126, 61, 240, 221, 178, 242, 159, 36, 138, 189, 0, 10, 125, 115, 167, 74, 81, 189, 67, 214, 106, 108, 209, 21, 222, 33, 144, 242, 174, 139, 72, 129, 68, 236, 199, 38, 88, 31, 229, 90, 120, 35, 177, 141, 167, 233, 16, 212, 6, 207, 101, 102, 40, 96, 51, 181, 73, 103, 162, 232, 49, 191, 86, 135, 33, 157, 60, 192, 105, 223, 40, 184, 171, 105, 83, 119, 95, 170, 137, 231, 56, 200, 17, 197, 58, 43, 23, 163, 56, 232, 216, 191, 84, 131, 102, 111, 112, 119, 108, 72, 13, 40, 234, 220, 237, 55, 158, 150, 246, 43, 198, 26, 247, 56, 192, 73, 149, 95, 173, 223, 174, 232, 118, 174, 112, 245, 168, 233, 76, 23, 157, 206, 11, 238, 3, 69, 242, 244, 210, 16, 85, 239, 136, 189, 224, 148, 231, 171, 105, 113, 47, 56, 63, 225, 58, 49, 227, 84, 123, 163, 39, 101, 116, 128, 70, 213, 93, 149, 246, 162, 200, 244, 173, 10, 209, 153, 192, 194, 119, 162, 197, 241, 228, 55, 193, 125, 47, 247, 72, 43, 85, 206, 108, 65, 87, 33, 245, 225, 35, 189, 88, 66, 157, 17, 134, 144, 91, 122, 39, 54, 35, 0, 158, 173, 212, 22, 157, 49, 104, 223, 122, 8, 24, 146, 147, 228, 62, 242, 181, 3, 142, 26, 178, 212, 158, 152, 107, 180, 10, 100, 71, 233, 4, 148, 108, 243, 166, 82, 218, 14, 127, 94, 165, 71, 4, 18, 3, 217, 182, 206, 250, 94, 17, 229, 26, 35, 104, 238, 117, 125, 0, 200, 108, 78, 240, 11, 250, 1, 76, 59, 57, 235, 116, 93, 11, 158, 195, 127, 36, 115, 59, 33, 0, 5, 144, 179, 56, 64, 61, 105, 173, 143, 227, 145, 196, 204, 87, 118, 168, 12, 13, 43, 107, 227, 185, 144, 94, 198, 31, 4, 210, 144, 228, 160, 184, 33, 167, 211, 35, 246, 151, 203, 77, 85, 130, 47, 118, 119, 203, 29, 180, 147, 131, 129, 102, 65, 56, 147, 36, 183, 101, 80, 64, 21, 24, 99, 214, 137, 22, 164, 170, 30, 233, 154, 67, 24, 27, 63, 138, 132, 149, 130, 101, 97, 86, 8, 199, 153, 18, 109, 166, 216, 190, 111, 128};
    logic [1:0] poly_ter [PARAM_N-1:0] = {0, 1, 3, 3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 1, 0, 1, 3, 0, 1, 0, 0, 0, 0, 1, 0, 0, 3, 0, 0, 0, 3, 0, 3, 0, 1, 3, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 3, 1, 3, 3, 0, 1, 0, 3, 0, 3, 0, 0, 3, 1, 1, 0, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 1, 3, 3, 0, 3, 3, 0, 3, 0, 1, 0, 0, 0, 1, 3, 0, 3, 0, 3, 3, 1, 3, 0, 3, 0, 0, 3, 3, 1, 3, 3, 1, 3, 3, 0, 3, 1, 1, 0, 1, 3, 1, 3, 1, 0, 3, 1, 3, 3, 1, 0, 0, 1, 1, 1, 0, 3, 3, 0, 1, 3, 3, 3, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 3, 0, 0, 0, 0, 3, 0, 1, 0, 3, 0, 3, 0, 0, 1, 3, 1, 3, 1, 3, 0, 0, 3, 3, 3, 0, 0, 1, 1, 0, 3, 1, 1, 3, 0, 0, 0, 0, 3, 0, 0, 1, 3, 3, 3, 0, 1, 1, 0, 0, 0, 0, 0, 3, 1, 0, 0, 3, 0, 3, 0, 3, 0, 0, 1, 1, 3, 1, 0, 3, 0, 0, 1, 0, 0, 1, 3, 0, 3, 0, 1, 1, 0, 1, 1, 0, 1, 0, 3, 0, 3, 0, 3, 3, 0, 3, 3, 0, 3, 1, 0, 0, 0, 3, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 0, 1, 0, 0, 0, 0, 1, 3, 1, 3, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 1, 1, 1, 0, 0, 0, 3, 1, 1, 0, 1, 1, 0, 3, 3, 0, 0, 3, 0, 3, 1, 3, 0, 0, 0, 1, 1, 3, 3, 0, 1, 3, 0, 0, 1, 3, 3, 0, 3, 3, 0, 0, 3, 0, 0, 0, 0, 0, 3, 1, 1, 1, 0, 0, 3, 3, 1, 0, 0, 3, 3, 0, 0, 3, 3, 0, 0, 3, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 3, 3, 0, 1, 1, 1, 0, 3, 3, 1, 0, 0, 3, 0, 0, 0, 0, 1, 1, 3, 1, 3, 0, 3, 0, 0, 0, 1, 3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 3, 0, 3, 1, 0, 0, 1, 3, 1, 1, 3, 0, 1, 0, 0, 3, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 3, 0, 3, 0, 3, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 0, 0, 0, 3, 0, 3, 0, 1, 0, 0, 3, 1, 3, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 1, 0, 3, 0, 1, 0, 3, 0, 0};
    
    initial
    begin
        #(`REF_CLK_PERIOD/2);
        clk = 1'b1;
        forever clk = #(`REF_CLK_PERIOD/2) ~clk;
    end
    
    initial
    begin
        rst = 0;
        enable_calc = 0;
        enable_write = 1;
        for (int i=0; i<510; i=i+5) begin
            in_1 = {poly_ter[i+2], poly_gen[i+2], poly_ter[i+1], poly_gen[i+1], poly_ter[i], poly_gen[i]};
            in_2 = {i, poly_ter[i+4], poly_gen[i+4], poly_ter[i+3], poly_gen[i+3]};
            #(`REF_CLK_PERIOD);
        end
        in_1 = {poly_ter[511], poly_gen[511],poly_ter[510], poly_gen[510]};
        in_2 = {12'h1FE, 20'b00000000000000000000};
        #(`REF_CLK_PERIOD);
        enable_write = 0;
        enable_calc = 1;
        #(`REF_CLK_PERIOD);
        #(`REF_CLK_PERIOD);
        wait (ready == 1'b1);
        enable_read = 1;
        #(`REF_CLK_PERIOD);
        in_1 = 0;
        for (int i=0; i<512; i=i+4) begin
            in_1 = i;
            #(`REF_CLK_PERIOD);
        end
        
    end
  
  mul_ternary_top mul_ternary_top_dut
  (
      .clk(clk),
      .rst(rst),
      .enable_write(enable_write),
      .enable_calc(enable_calc),
      .enable_read(enable_read),
      .in_1(in_1),
      .in_2(in_2),
      .out_1(out_1),
      .ready(ready)
  );
    
endmodule
