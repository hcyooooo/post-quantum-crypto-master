`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Technical University of Munich
// Engineer: Tim Fritzmann
// 
// Create Date: 01/27/2020
// Module Name: cal_syndrome_tb
// Project Name: Post-Quantum Cryptography
// 
//////////////////////////////////////////////////////////////////////////////////


`define CLK_PERIOD       40.00ns      // 25 MHz

module cal_syndrome_tb;
//    parameter PARAM_M = 4;
//    parameter PARAM_ALPHA = 1;
    parameter PARAM_M = 9;
    parameter PARAM_ALPHA = 4;
//    parameter PARAM_ECC_BITS = 171;
//    parameter PARAM_ECC_BITS = 171;
    parameter PARAM_ECC_BITS = 160;
    parameter PARAM_LOG_ECC_BITS = 8;
    logic clk;
    logic rst;    
    logic [PARAM_ECC_BITS-1:0] in_1;
    logic [PARAM_M-1:0] out_1;


    cal_syndrome #(.PARAM_M(PARAM_M), .PARAM_ALPHA(PARAM_ALPHA), .PARAM_ECC_BITS(PARAM_ECC_BITS), .PARAM_LOG_ECC_BITS(PARAM_LOG_ECC_BITS)) mul_general_dut
    (
        .clk(clk),
        .rst(rst),    
        .in_1(in_1),
        .out_1(out_1)
    );
    
    initial
    begin
//       in_1 = 4'b1111;
//       in_2 = 4'b0100;
//       in_1 = 171'b000000000000110110010010011000001100101010110100001001101100000100001001111100100101110011000011100101111100111010000110111111000000011111001000100101110100101110011110011;
//       in_1 = 192'b111101100110000000000000000000000110110010010011000001100101010110100001001101100000100001001111100100101110011000011100101111100111010000110111111000000011111001000100101110100101110011110011;
//         in_1 = 171'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
//         in_1 = 171'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111;
//       in_1 = 171'b110011110011101001011101001000100111110000000111111011000010111001111101001110000110011101001001111100100001000001101100100001011010101001100000110010010011011000000000000;
//       in_1 = 0;
//       in_1 = 144'b0000000000000000011011001010001110001110101110100010011111110001000110100110011101110010110100011010100111001101011100101110011001011101011001111001000110111100;
//       in_1 = 164'b0011110110001001111001101011101001100111010011101011001110010101100010110100111011100110010110001000111111100100010111010111000111000101001101100000000000000000;
       in_1 = 160'b0011110110001001111001101011101001100111010011101011001110010101100010110100111011100110010110001000111111100100010111010111000111000101001101100000000000000000;
       in_1 = 160'b0000000000000000011011001010001110001110101110100010011111110001000110100110011101110010110100011010100111001101011100101110011001011101011001111001000110111100;
       rst = 0;
       #(`CLK_PERIOD);
       rst = 1;
       #(`CLK_PERIOD*2);
       rst = 0;
       
       
    end
    
    initial
    begin
      clk = 1'b0;
      #(`CLK_PERIOD/2);
      clk = 1'b1;
      forever clk = #(`CLK_PERIOD/2) ~clk;
    end
       

endmodule

